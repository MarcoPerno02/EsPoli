** dsd
V1 1 0 dc 3
R1 1 0 1
R2 2 1 1.5
E1 3 2 1 2 2
R4 3 0 3
.op
.end
