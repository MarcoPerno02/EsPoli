*www
R9 1 0 22000
Rid 1 2 1000000
R8 2 0 10000
R10 1 3 100000
Ro 3 4 100
E1 4 0 2 1 200000
VP 3 0 400
.op
.end
