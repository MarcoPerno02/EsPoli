*www
VP 1 0 400
Rid 1 2 1000000
R2 2 0 12000
Routand1 3 2 100100
E1 3 0 1 2 200000
.op
.end
