*ssa
I1 0 1 1
R1 1 0 2
R2 1 2 8
G1 2 0 1 0 2
R3 2 3 5
Vp 3 0 4
.op
.end
