* cicuito da analizzare epr la scimmia
v1 2 0 dc 5
r3 2 0 10k
e 3 0 2 1 999k
r1 3 1 20k
r2 1 0 10k
.op
.end
