*www
VP 1 0 600
R9 2 1 22000
Rid 2 3 1000000
R8 3 0 10000
R10 2 4 100000
Ro 4 5 100
E1 5 0 3 2 200000
.op
.end
