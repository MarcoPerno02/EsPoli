*aa
R1 2 3 3
Vd 3 0 dc 0
Vs 2 0 dc -1
F1 1 0 Vd 3
Is 2 1 1
R2 1 0 3
Vp 1 0 dc 1
.op
.end
