*** e
V1 2 0 8
R1 1 2 6
Vd 1 2 0
I1 1 0 2
R2 1 4 3
H2 4 0 Vd 3
.op
.end
