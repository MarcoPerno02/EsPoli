**aaaa
R1 0 2 3
R2 0 1 2
I1 0 1 3
E1 1 2 0 1 1
R3 0 1 2
.op
.end
