*www
Rid 0 2 1000000
R2 2 0 12000
Rout 3 4 100000
R1 4 2 100
E1 3 0 0 2 200000
VP 4 0 300
.op
.end
