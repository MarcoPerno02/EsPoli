*www
V1 3 0 1
R4 3 1 2
R3 1 0 6
R2 1 2 2
R1 2 0 4
E1 1 2 2 0 2
.op
.end
