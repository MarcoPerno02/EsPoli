E1;
Vg 1 0 100;
R1 1 2 250
R2 2 0 750
.op
.end
