*aaaa
v1 1 0 dc 10
r1 1 2 3k
r2 0 2 2k
r3 0 3 10k
r4 3 4 20k
r5 0 4 2k
XOA1 2 3 4 opamp

.SUBCKT OPAMP 1 2 3
E0A 3 0 1 2 1e8
.ENDS

.op
.end



